,id,title,release_date,overview,popularity,vote_average
0,533514,Violet Evergarden: The Movie,2020-09-18,"As the world moves on from the war and technological advances bring changes to her life, Violet still hopes to see her lost commanding officer again.",7.412,8.3
1,975,Paths of Glory,1957-10-25,A commanding officer defends three scapegoats on trial for a failed offensive that occurred within the French Army in 1916.,6.382,8.259
2,637920,Miracle in Cell No. 7,2019-10-10,"Separated from his daughter, a father with an intellectual disability must prove his innocence when he is jailed for the death of a commander's child.",7.17,8.3
3,10376,The Legend of 1900,1998-10-28,"The story of a virtuoso piano player who lives his entire life aboard an ocean liner. Born and raised on the ship, 1900 (Tim Roth) learned about the outside world through interactions with passengers, never setting foot on land, even for the love of his life. Years later, the ship may be destroyed, and a former band member fears that 1900 may still be aboard, willing to go down with the ship.",4.91,8.3
4,8587,The Lion King,1994-06-15,"Young lion prince Simba, eager to one day become king of the Pride Lands, grows up under the watchful eye of his father Mufasa; all the while his villainous uncle Scar conspires to take the throne for himself. Amid betrayal and tragedy, Simba must confront his past and find his rightful place in the Circle of Life.",36.209,8.255
5,29259,Le Trou,1960-03-18,"Four prison inmates have been hatching a plan to literally dig out of jail when another prisoner, Claude Gaspard, is moved into their cell. They take a risk and share their plan with the newcomer. Over the course of three days, the prisoners and friends break through the concrete floor using a bed post and begin to make their way through the sewer system -- yet their escape is anything but assured.",4.475,8.3
6,670,Oldboy,2003-11-21,"With no clue how he came to be imprisoned, drugged and tortured for 15 years, a desperate man seeks revenge on his captors.",18.301,8.253
7,630566,Clouds,2020-10-09,"Young musician Zach Sobiech discovers his cancer has spread, leaving him just a few months to live. With limited time, he follows his dream and makes an album, unaware that it will soon be a viral music phenomenon.",4.893,8.2
8,572154,Rascal Does Not Dream of a Dreaming Girl,2019-06-15,"In Fujisawa, Sakuta Azusagawa is in his second year of high school. Blissful days with his girlfriend and upperclassman, Mai Sakurajima, are interrupted by the appearance of his first crush, Shoko Makinohara.",5.267,8.246
9,1160164,TAYLOR SWIFT | THE ERAS TOUR,2023-10-13,"The cultural phenomenon continues on the big screen! Immerse yourself in this once-in-a-lifetime concert film experience with a breathtaking, cinematic view of the history-making tour.",8.186,8.2
10,995133,"The Boy, the Mole, the Fox and the Horse",2022-12-25,"The unlikely friendship of a boy, a mole, a fox and a horse traveling together in the boy's search for home.",7.217,8.245
11,447362,Life in a Year,2020-11-27,"A 17 year old finds out that his girlfriend is dying, so he sets out to give her an entire life, in the last year she has left.",8.648,8.245
12,508965,Klaus,2019-11-08,"When Jesper distinguishes himself as the Postal Academy's worst student, he is sent to Smeerensburg, a small village located on an icy island above the Arctic Circle, where grumpy inhabitants barely exchange words, let alone letters. Jesper is about to give up and abandon his duty as a postman when he meets local teacher Alva and Klaus, a mysterious carpenter who lives alone in a cabin full of handmade toys.",7.556,8.243
13,527641,Five Feet Apart,2019-03-14,"Seventeen-year-old Stella spends most of her time in the hospital as a cystic fibrosis patient. Her life is full of routines, boundaries and self-control — all of which get put to the test when she meets Will, an impossibly charming teen who has the same illness. There's an instant flirtation, though restrictions dictate that they must maintain a safe distance between them. As their connection intensifies, so does the temptation to throw the rules out the window and embrace that attraction.",12.904,8.241
14,504253,I Want to Eat Your Pancreas,2018-09-01,"After his classmate and crush is diagnosed with a pancreatic disease, an average high schooler sets out to make the most of her final days.",7.285,8.2
15,299534,Avengers: Endgame,2019-04-24,"After the devastating events of Avengers: Infinity War, the universe is in ruins due to the efforts of the Mad Titan, Thanos. With the help of remaining allies, the Avengers must assemble once more in order to undo Thanos' actions and restore order to the universe once and for all, no matter what consequences may be in store.",30.301,8.24
16,25237,Come and See,1985-10-17,"The invasion of a village in Byelorussia by German forces sends young Florya into the forest to join the weary Resistance fighters, against his family's wishes. There he meets a girl, Glasha, who accompanies him back to his village. On returning home, Florya finds his family and fellow peasants massacred. His continued survival amidst the brutal debris of war becomes increasingly nightmarish, a battle between despair and hope.",8.456,8.2
17,299536,Avengers: Infinity War,2018-04-25,"As the Avengers and their allies have continued to protect the world from threats too large for any one hero to handle, a new danger has emerged from the cosmic shadows: Thanos. A despot of intergalactic infamy, his goal is to collect all six Infinity Stones, artifacts of unimaginable power, and use them to inflict his twisted will on all of reality. Everything the Avengers have fought for has led up to this moment - the fate of Earth and existence itself has never been more uncertain.",64.75,8.237
18,490132,Green Book,2018-11-16,"Tony Lip, a bouncer in 1962, is hired to drive pianist Don Shirley on a tour through the Deep South in the days when African Americans, forced to find alternate accommodations and services due to segregation laws below the Mason-Dixon Line, relied on a guide called The Negro Motorist Green Book.",24.938,8.2
19,265177,Mommy,2014-09-19,"A peculiar neighbor offers hope to a recent widow who is struggling to raise a teenager who is unpredictable and, sometimes, violent.",5.214,8.2
